package ArmFilePaths is 

	--	Pfad zum Testvektorverzeichnis, betriebssystem- und und Projektabhängig;
	constant TESTVECTOR_FOLDER_PATH : STRING := "/home/tu-berlin.de/azizlazzem/irb-ubuntu/Desktop/HWPTI/VECTORS/";

end package ArmFilePaths;

package body ArmFilePaths is
end package body ArmFilePaths;
